module mod1();

mod3 mod3_inst1();


endmodule