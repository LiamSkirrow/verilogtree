module mod2();

mod1 mod1_inst1();


endmodule