module 
    mod4();



endmodule
