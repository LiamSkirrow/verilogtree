module mod3();




endmodule