module mod0 ();


mod3 mod3_inst0();
mod1 mod1_instAnother();


endmodule
