   module    mod1 ();

mod3 mod3_inst1();

// comment with word module in it

// module comment0 (


endmodule

/* 
// module comment1 (

*/
