module altTop();


mod2 mod2_instX();


endmodule
