module altTop();


mod3 mod3_instX();


endmodule