module mod0();


mod3 mod3_inst0();


endmodule