module
    mod3
();

mod4 mod4_inst();


endmodule
